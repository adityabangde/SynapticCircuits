.title RC_Low_Pass_Filter

frequency domain
.end

